module and_gate(input a,b,output out1);
  assign out1= a & b;
endmodule
module and_gate1(input x,y,z,output out2);
  assign out2 = x & y & z;
endmodule
