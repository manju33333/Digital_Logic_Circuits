// Code your design here
module exor_gate(input a,b,output out);
  assign out = a ^ b;
endmodule