module half_subtractor_tb;
reg A, B;
wire Diff, Borrow;

half_subtractor uut (.A(A), .B(B), .Diff(Diff), .Borrow(Borrow));

initial begin
    A=0; B=0; #10;
    A=0; B=1; #10;
    A=1; B=0; #10;
    A=1; B=1; #10;
    $finish;
end
endmodule
