// Code your design here
module exnor_gate(input a,b,output out);
  assign out = a ~^ b;
endmodule